entity testbench is
end entity;
