library ieee;
use ieee.std_logic_1164.all;

entity clock is
end entity;

architecture clock_arch of clock is
begin
end architecture;