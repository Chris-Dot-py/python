library ieee;
use ieee.std_logic_1164.all;

entity tb_clock is
end entity;

architecture tb_clock_arch of tb_clock is
begin
end architecture;