library ieee;
use ieee.std_logic_1164.all;

entity testfile is
end entity;

architecture testfile_arch of testfile is
begin
end architecture;